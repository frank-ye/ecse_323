library verilog;
use verilog.vl_types.all;
entity gA8_comp7_vlg_vec_tst is
end gA8_comp7_vlg_vec_tst;
