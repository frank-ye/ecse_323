library verilog;
use verilog.vl_types.all;
entity g08_rules_vlg_check_tst is
    port(
        legal_play      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g08_rules_vlg_check_tst;
