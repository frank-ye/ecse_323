library verilog;
use verilog.vl_types.all;
entity g08_adder_vlg_vec_tst is
end g08_adder_vlg_vec_tst;
