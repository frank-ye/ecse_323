library verilog;
use verilog.vl_types.all;
entity DIVIDE10_vlg_vec_tst is
end DIVIDE10_vlg_vec_tst;
