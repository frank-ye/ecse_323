library verilog;
use verilog.vl_types.all;
entity g08_pulseGenerator_vlg_vec_tst is
end g08_pulseGenerator_vlg_vec_tst;
