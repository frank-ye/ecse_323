library verilog;
use verilog.vl_types.all;
entity TIME13_vlg_vec_tst is
end TIME13_vlg_vec_tst;
