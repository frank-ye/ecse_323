library verilog;
use verilog.vl_types.all;
entity gA8_lab1_vlg_vec_tst is
end gA8_lab1_vlg_vec_tst;
