library verilog;
use verilog.vl_types.all;
entity FLOOR13_vlg_vec_tst is
end FLOOR13_vlg_vec_tst;
