library verilog;
use verilog.vl_types.all;
entity test_bed_vlg_vec_tst is
end test_bed_vlg_vec_tst;
