library verilog;
use verilog.vl_types.all;
entity gA8_lab1_vlg_check_tst is
    port(
        AeqB            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end gA8_lab1_vlg_check_tst;
